
class scoreboard;


function new(); // Get register values and fetched instruction pc etc here
begin
    
end


endclass

