package alu_pkg;

	`include "mips_16_defs.v"
	`include "alu_defs.sv"

	`include "transaction.sv"
	`include "alu_scoreboard.sv"
	`include "alu_driver.sv"
	`include "alu_monitor.sv"
	`include "alu_coverage.sv"


endpackage : alu_pkg