
package hd_pkg;

	`include "mips_16_defs.v"
	`include "hd_defs.sv"

	`include "transaction.sv"
	`include "hd_scoreboard.sv"
	`include "hd_driver.sv"
	`include "hd_monitor.sv"
	`include "hd_coverage.sv"


endpackage : hd_pkg